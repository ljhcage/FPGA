/***************************************************************************************
FILE NAME      :     Frequency_Counter
AUTHOR         :     Crazy Bingo
FUNCTION       :     MCU430 and CPLD to control the Frequency counter 
FEATURE        :     EPM240T100C5N
SETUP TIME     :     2010/5/6
***************************************************************************************/
module Frequency_Counter(
						input				CLOCK_50,		//����ʱ��
						input				RST_n,		//ϵͳ��λ�����ź�	
						
						input				Fx,			//�����ź�Ƶ��	
						//��Fx�����ؼ�⣬ʵ����Fx������ͬ�����Ӷ���֤������2�Ա����źŸպ�Ϊ����������,0���
						input				Cnt_Sel,	//Ƶ�ʼ���ѡ��cnt_Fb,cnt_Fx��
						input		[1:0]	Byte_Sel,	//CLK��������ַλѡ				
						
						output	reg			Finish,		//The Measure of the frequency is finished 		
						output	reg	[7:0]	Freq_Data	//����Ƶ�ʼ�
						);	
													//999_999999=27'h3b9ac9ff
reg			cnt_EN;		//�������ſ����źţ�ͨ��D��������ʱ�Ӵﵽͬ
reg			Finish_r;
reg	[31:0]	cnt_Fb;		//��׼Դ	Fb 	������	//32'hFFFFFFFF=32'd4294967295=429 MHz
reg	[31:0]	cnt_Fx;		//�����ź�	Fx	������
reg	[26:0]	cnt_1s;		
reg			cnt_Flag;
reg	[15:0]	cnt;


always@(posedge CLOCK_50 or negedge RST_n)
begin
	if(!RST_n)
		begin
		cnt_1s <= 0;
		cnt_Flag <= 0;
		Finish_r <= 0;
		end
	else
		begin
		if(cnt_1s < 27'd50_000000)	//2s
			begin
			cnt_1s <= cnt_1s+1'b1;
			cnt_Flag <= 1;
			Finish_r <= 0;
			end
		else
			begin
			cnt_1s <= cnt_1s;
			cnt_Flag <= 0;		//The signal means that it has reach the time of 1S
			Finish_r <= 1;		//Lock the signal Finish for math calculation
			end
		end
end

//�Ⱦ���Ƶ�ʼ��ſ����ź�
//Gate�Ŀ��Tc�ͷ�����ʱ�䶼����ֱ��Ӱ�����ʹ���ź�EN��EN�����ڱ����ź�fx�����ظı䣬
//�Ӷ���֤�˱����źű�������������������������nTx�����뱻���źŵ�Ƶ���޹�
always@(posedge Fx or negedge RST_n)	//D������ʵ�ֶԱ����ź�fx�����ؼ�⣬ʵ���ſ��ź���fx������ͬ����
begin									//�Ӷ���֤������2�Ա����źż����պ�Ϊ���������ڣ�����
	if(!RST_n)
		begin
		cnt_EN <= 0;
		Finish <= 0;
		end
	else								//�ڱ����ź�fb�����ص���t2ʱ��D������Q�˲ű���1
		begin
		if(cnt_Flag==1'b1)
			cnt_EN <= 1;				//ʹ������1�ͼ�����2��ENͬʱΪ1����������ʼ������ϵͳ��������������ڡ�
		else
			cnt_EN <= 0;
		
		if(Finish_r==1'b1)
			Finish <= 1;
		else
			Finish <= 0;
		end
end

////Fb ��׼Դ����ģ��
always@(posedge CLOCK_50 or negedge RST_n)		
begin
	if(!RST_n)
		cnt_Fb <= 0;
	else
		begin
		if(cnt_Flag==1'b1)//if(EN==1'b1)
			cnt_Fb <= cnt_Fb+1'b1;
		else
			cnt_Fb <= cnt_Fb;	//Locked		
		end
end
//
////FX �����źż���ģ��
always@(posedge Fx  or negedge RST_n)		
begin
	if(!RST_n)
		cnt_Fx <= 0;
	else
		begin
		if(cnt_Flag==1'b1)//if(EN==1'b1)
			cnt_Fx <= cnt_Fx+1'b1;
		else
			cnt_Fx <= cnt_Fx;	//Locked		
		end
end

//cnt_Fb,cnt_Fb		32λ���������ֳ�2��16λ�ͳ�
//Freq_Data[15:0]	16λ��������
//MCU  				�������ݲ�����Ӧ����
//always@(RD,Cnt_Sel,Byte_Sel,cnt_Fb,cnt_Fx)

//always@(posedge CLOCK_50 or negedge RST_n)
always@(Cnt_Sel,Byte_Sel,cnt_Fb,cnt_Fx)
begin
//	cnt_Fb=32'd50_000000;	//32'h02_FA_F0_80
	//cnt_Fx=32'd1000000;	   //32'h00_98_96_80
	case({Cnt_Sel,Byte_Sel})
	4'b000	:		Freq_Data <= cnt_Fb[7:0];	//Fb ��׼Դ����ģ��
	4'b001	:		Freq_Data <= cnt_Fb[15:8];
	4'b010	:		Freq_Data <= cnt_Fb[23:16];
	4'b011	:		Freq_Data <= cnt_Fb[31:24];	
	4'b100	:		Freq_Data <= cnt_Fx[7:0];	//Fx �����źż���ģ��
	4'b101	:		Freq_Data <= cnt_Fx[15:8];
	4'b110	:		Freq_Data <= cnt_Fx[23:16];
	4'b111	:		Freq_Data <= cnt_Fx[31:24];
	endcase 	
end

endmodule
